`include "./src/alu.v"
`include "./src/control_unit.v"
`include "./src/mux.v"
`include "./src/memory.v"
`include "./src/register_file.v"
`include "./src/alu_control.v"
`include "./src/inst_mem.v"
`include "./src/pc.v"

module cpu(
    input clk,
    input rst,
);




endmodule